`timescale 1ns/1ps
module TimeController(
  
);

endmodule // TimeController