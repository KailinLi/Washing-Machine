`timescale 1ns/1ps
module View(
  
);

endmodule // View